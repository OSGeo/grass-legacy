src/libes/vask
src/libes/segment
src/libes/rowio
src/libes/raster
src/libes/lock
src/libes/imagery
src/libes/icon
src/libes/gis
src/libes/dlg
src/libes.datetime
src/libes/dbmi
src/libes/geom
src/libes/proj
src/libes/display
src/libes/dig_atts
src/libes/coorcnv
src/libes/btree
src/libes/ibtree
src/libes/linkm
src/libes/bitmap
src/libes/D
src/mapdev/libes
src/mapdev/Vlib
src/mapdev/diglib
src/display/devices/lib
src/display/devices/monitorcap
src/fonts/for_grass
src/front.end
src/display/d.3d
src/display/d.ask
src/display/d.colormode
src/display/d.colors
src/display/d.colortable
src/display/d.display
src/display/d.erase
src/display/d.font
src/display/d.frame
src/display/d.geodesic
src/display/d.graph
src/display/d.grid
src/display/d.his
src/display/d.histogram
src/display/d.icons
src/display/d.label
src/display/d.legend
src/display/d.mapgraph
src/display/d.measure
src/display/d.menu
src/display/d.mon
src/display/d.mouse
src/display/d.p.labels
src/display/d.points
src/display/d.profile
src/display/d.rast
src/display/d.rgb
src/display/d.rhumbline
src/display/d.save
src/display/d.scale
src/display/d.sites
src/display/d.text
src/display/d.title
src/display/d.vect
src/display/d.what.rast
src/display/d.what.vect
src/display/d.where
src/display/d.zoom
src/imagery/i.ask
src/imagery/i.cca
src/imagery/i.class
src/imagery/i.colors
src/imagery/i.composite
src/imagery/i.fft
src/imagery/i.find
src/imagery/i.grey.scale
src/imagery/i.group
src/imagery/i.maxlik
src/imagery/i.pca
src/imagery/i.points
src/imagery/i.rectify
src/imagery/i.rgb.his
src/imagery/i.tape.mss
src/imagery/i.tape.mss.h
src/imagery/i.tape.other
src/imagery/i.tape.tm
src/imagery/i.target
src/imagery/i.zc
src/general/g.access
src/general/g.ask
src/general/g.filename
src/general/g.findfile
src/general/g.gisenv
src/general/g.help
src/general/g.manual
src/general/g.mapsets
src/general/g.region
src/general/g.tempfile
src/general/g.setproj
src/general/g.version
src/general/gis
src/general/manage
src/mapdev/v.area
src/mapdev/v.build
src/mapdev/v.cadlabel
src/mapdev/v.clean
src/mapdev/v.digit
src/mapdev/v.from.3
src/mapdev/v.import
src/mapdev/v.in.ascii
src/mapdev/v.in.dlg
src/mapdev/v.in.dxf
src/mapdev/v.mkgrid
src/mapdev/v.mkquads
src/mapdev/v.out.dlg
src/mapdev/v.out.dxf
src/mapdev/v.patch
src/mapdev/v.prune
src/mapdev/v.spag
src/mapdev/v.stats
src/mapdev/v.support
src/mapdev/v.to.rast
src/mapdev/v.transform
src/mapdev/v.trim
src/mapdev/georef
src/paint/Interface
src/paint/Drivers
src/paint/Drivers/NULL
src/paint/Drivers/act2
src/paint/Drivers/diablo.c150
src/paint/Drivers/epson.lq2500
src/paint/Drivers/genicom3310
src/paint/Drivers/ppm
src/paint/Drivers/preview
src/paint/Drivers/preview2
src/paint/Drivers/shinko635
src/paint/Drivers/tek4695
src/paint/Drivers/tek4697
src/paint/Drivers/versatec/driver
src/paint/Drivers/versatec/3236
src/paint/Drivers/versatec/3236.fast
src/paint/Drivers/versatec/3236.slow
src/paint/Drivers/xerox4020
src/paint/Programs
src/paint/Tests
src/raster/r.average
src/raster/r.basins.fill
src/raster/r.binfer
src/raster/r.buffer
src/raster/r.cats
src/raster/r.clump
src/raster/r.coin
src/raster/r.colors
src/raster/r.combine
src/raster/r.compress
src/raster/r.covar
src/raster/r.cross
src/raster/r.describe
src/raster/r.drain
src/raster/r.grow
src/raster/r.in.ascii
src/raster/r.in.ll
src/raster/r.infer
src/raster/r.info
src/raster/r.kappa
src/raster/r.los
src/raster/r.mapcalc
src/raster/r.mfilter
src/raster/r.neighbors
src/raster/r.null
src/raster/r.out.ascii
src/raster/r.patch
src/raster/r.poly
src/raster/r.profile
src/raster/r.quant
src/raster/r.random
src/raster/r.reclass
src/raster/r.recode
src/raster/r.report
src/raster/r.resample
src/raster/r.rescale
src/raster/r.slope.aspect
src/raster/r.stats
src/raster/r.support
src/raster/r.surf.idw
src/raster/r.surf.idw2
src/raster/r.transect
src/raster/r.volume
src/raster/r.watershed
src/raster/r.weight
src/raster/r.what
src/sites/s.in.ascii
src/sites/s.menu
src/sites/s.out.ascii
src/sites/s.surf.idw
src/sites/s.to.rast
src/sites/sroff
src/misc/m.dem.examine
src/misc/m.dmaUSGSread
src/misc/m.dted.examine
src/misc/m.dted.extract
src/misc/m.examine.tape
src/misc/m.gc2ll
src/misc/m.ll2gc
src/misc/m.ll2u
src/misc/m.region.ll
src/misc/m.rot90
src/misc/m.u2ll
src/scripts
src/display/d.labels
src/display/d.rast.arrow
src/display/d.rast.edit
src/display/d.rast.num
src/display/d.rast.zoom
src/imagery/i.cluster
src/imagery/i.gensig
src/imagery/i.gensigset
src/imagery/i.in.erdas
src/imagery/i.ortho.photo
src/imagery/i.quantize
src/imagery/i.rectify2
src/imagery/i.smap
src/imagery/i.tape.spot
src/imagery/i.tape.tm.fast
src/imagery/i.vpoints
src/mapdev/moss
src/mapdev/v.alabel
src/mapdev/v.apply.census
src/mapdev/v.cutter
src/mapdev/v.in.arc
src/mapdev/v.in.tig.basic
src/mapdev/v.in.tig.lndmk
src/mapdev/v.in.transects
src/mapdev/v.out.arc
src/mapdev/v.proj
src/mapdev/v.reclass
src/mapdev/v.to.sites
src/paint/Programs/p.map.new/cmd
src/ps.map
src/raster/r.colors.paint
src/raster/r.contour
src/raster/r.cost
src/raster/r.digit
src/raster/r.in.poly
src/raster/r.in.sunrast
src/raster/r.line
src/raster/r.mask.points
src/raster/r.median
src/raster/r.mode
src/raster/r.out.tga
src/raster/r.rescale.eq
src/raster/r.surf.contour
src/raster/r.surf.contour/cmd
src/raster/r.thin
src/raster/r.weight2
src/sites/s.surf.tps
src/misc/m.dem.extract
src/misc/m.flip
src/misc/m.in.pl94.db3
src/misc/m.in.stf1.db3
src/misc/m.in.stf1.tape
src/misc/m.lulc.USGS
src/misc/m.lulc.read
src/misc/m.proj
src/misc/m.tiger.region
#######################################
